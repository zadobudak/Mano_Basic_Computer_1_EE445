//Don't change the module I/O
module BC_I (
input clk,
input FGI,
output [11:0] PC,
output [11:0] AR,
output [15:0] IR,
output [15:0] AC,
output [15:0] DR
);

// Instantiate your datapath and controller here, then connect them.

endmodule